module fpga_top;
    reg a;
    wire b;
    two _two(a, b);
endmodule
