module fpga_top;
endmodule
